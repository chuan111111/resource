module lab31 (
    input [1:0] a,b,c,d,
    
    output [2:0] sum
    
);
assign sum[0]=~a[1]&~a[0]&~b[1]&b[0]|~a[0]&~a[1]&b[0]&b[1]|~a[1]&a[0]&~b[1]&~b[0]|~a[1]&a[0]&b[1]&~b[0]|a[1]&~a[0]&~b[1]&b[0]|a[1]&~a[0]&b[1]&b[0]|a[1]&a[0]&~b[1]&~b[0]|a[1]&a[0]&b[1]&~b[0];
assign  sum[1]=~a[1]&~a[0]&b[1]&~b[0]|~a[1]&~a[0]&b[1]&b[0]|~a[1]&a[0]&~b[1]&b[0]|~a[1]&a[0]&b[1]&~b[0]|a[1]&~a[0]&~b[1]&~b[0]|a[1]&~a[0]&~b[1]&b[0]|a[1]&a[0]&~b[1]&~b[0]|a[1]&a[0]&b[1]&b[0];
assign  sum[2]=~a[1]&a[0]&b[1]&b[0]|a[1]&~a[0]&b[1]&~b[0]|a[1]&~a[0]&b[1]&b[0]|a[1]&a[0]&~b[1]&b[0]|a[1]&a[0]&b[1]&~b[0]|a[1]&a[0]&b[1]&b[0];
assign sum[0]=sum[1]&sum[2];
    
endmodule