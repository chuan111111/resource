module lab4_sim ( );
    ports
);
    
endmodule