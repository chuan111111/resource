module lab32 (
    input  a,b,
    output  sum
);

assign sum=a+b;
  
endmodule