module lab4 (
    input x,
    input y,
    input z
);
assign
    
endmodule